module Adder4(input logic [31:0] adress,
						output logic [31:0] adressp4);
						
assign new_adress = adress + 32'b00000000000000000000000000000100;

endmodule
